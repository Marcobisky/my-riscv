LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity DIG_LUT_LUT_inst_Decoder is
  port (
    n0: in std_logic;
    n1: in std_logic;
    n2: in std_logic;
    n3: in std_logic;
    n4: in std_logic;
    n5: in std_logic;
    n6: in std_logic;

    p_out: out std_logic_vector (3 downto 0)
);
end DIG_LUT_LUT_inst_Decoder;

architecture Behavioral of DIG_LUT_LUT_inst_Decoder is
  type mem is array ( 0 to 127) of std_logic_vector (3 downto 0);
  constant my_lut : mem := (
    "0000", "0000", "0000", "0101", "0000", "0000", "0000", "0000", "0000", 
    "0000", "0000", "0000", "0000", "0000", "0000", "1011", "0000", "0000", 
    "0000", "0010", "0000", "0000", "0000", "1001", "0000", "0000", "0000", 
    "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1000", 
    "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", 
    "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0000", "0000", 
    "0000", "1010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", 
    "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", 
    "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", 
    "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", 
    "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", 
    "0001", "0000", "0000", "0000", "0100", "0000", "0000", "0000", "0000", 
    "0000", "0000", "0000", "0110", "0000", "0000", "0000", "0011", "0000", 
    "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", 
    "0000", "1111");
  signal temp : std_logic_vector(6 downto 0);
begin
  temp <= n6 & n5 & n4 & n3 & n2 & n1 & n0;
  p_out <= my_lut(to_integer(unsigned(temp)));
end Behavioral;